package master_package;
typedef enum {ERROR,OKAY}HRESP_E;
typedef enum {BYTE,HALF_WORD,WORD}HSIZE_E;
typedef enum {IDLE,BUSY,NONSEQ,SEQ}HTRANS_E;
typedef enum {SINGLE,INCR}HBURST_E;


endpackage
